`define R_TYPE_OP     7'b0110011
`define I_TYPE_ALU_OP 7'b0010011
`define LW_OP         7'b0000011
`define SW_OP         7'b0100011
`define BRANCH_OP     7'b1100011
`define JAL_OP        7'b1101111
`define JALR_OP       7'b1100111
`define LUI_OP        7'b0110111
`define AUIPC_OP     7'b0010111